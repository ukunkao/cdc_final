
module flip_flop_synch_1bit(
    input wire a_clk,            
    input wire a_rst_n,          
    input wire b_clk,           
    input wire b_rst_n,         
    input wire  async_data,   
    output reg  sync_data     
);


    reg  stage1;
    reg  stage2;


    always @(posedge a_clk or posedge a_rst_n) begin
        if (a_rst_n) begin
            stage1 <= 1'b0;
        end else begin
            stage1 <= async_data;
        end
    end

    always @(posedge b_clk or posedge b_rst_n) begin
        if (b_rst_n) begin
            stage2 <= 1'b0;
            sync_data <= 1'b0;
        end else begin
            stage2 <= stage1;  
            sync_data <= stage2;  
        end
    end
endmodule


